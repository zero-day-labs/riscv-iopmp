// Author: Luís Cunha
// Date: 23/02/2024
// Acknowledges: Manuel Rodríguez <manuel.cederog@gmail.com>
//
// Description: AXI4 Boundary Checker module for RISC-V IOPMP:
//              Checks whether an AXI transaction crosses a 4-kiB address boundary,
//              which is illegal in AXI4 transactions.

/* verilator lint_off WIDTH */

module rv_iopmp_axi4_bc (
    // AxVALID
    input  logic                    request_i,
    // AxADDR
    input  logic [64-1:0]           addr_i,
    // AxBURST
    input  axi_pkg::burst_t         burst_type_i,
    // AxLEN
    input  axi_pkg::len_t           burst_length_i,
    // AxSIZE
    input  axi_pkg::size_t          n_bytes_i,

    // To indicate valid requests or boundary violations
    output logic                    allow_request_o,
    output logic                    bound_violation_o,
    output logic [64-1:0]           wrap_boundary_o
);

always_comb begin : boundary_check

    allow_request_o   = 1'b0;
    bound_violation_o = 1'b0;
    wrap_boundary_o   = '0;

    // Request received
    if (request_i) begin

        // Consider burst type, N of beats and size of the beat (always 64 bits) to calculate number of bytes accessed:
        case (burst_type_i)

            // BURST_FIXED: The final address is Start Addr + 8 (ex: ARADDR + 8)
            axi_pkg::BURST_FIXED: begin
                // May be optimized with bitwise AND
                if (((addr_i & 12'hfff) + (1'b1 << n_bytes_i)) < (1'b1 << 12)) begin
                    allow_request_o   = 1'b1;     // Allow transaction
                end

                // Boundary violation
                else begin
                    bound_violation_o = 1'b1;
                end
            end

            // BURST_WRAP: The final address is the Wrap Boundary (Lower address) + size of the transfer
            axi_pkg::BURST_WRAP: begin
                // wrap_boundary = (start_address/(number_bytes*burst_length_i)) * (number_bytes*burst_length_i)
                // address_n = wrap_boundary + (number_bytes * burst_length_i)

                // by spec, N of transfers must be {2, 4, 8, 16}
                // So, ARLEN must be {1, 3, 7, 15}
                logic [2:0] log2_len;
                case (burst_length_i)
                    8'd1: log2_len = 3'b001;
                    8'd3: log2_len = 3'b010;
                    8'd7: log2_len = 3'b011;
                    8'd15: log2_len = 3'b100;
                    default: log2_len = 3'b111;  // invalid
                endcase

                // As we need this, no need to replicate this logic elsewhere
                // The lowest address within a wrapping burst
                // Wrap_Boundary = (INT(Start_Address / (Burst_Length x Number_Bytes))) x (Burst_Length x Number_Bytes)
                wrap_boundary_o = (addr_i >> (log2_len + n_bytes_i)) << (log2_len + n_bytes_i);

                // Check if the highest address crosses a 4 kiB boundary (Highest Addr - Lower Addr >= 4kiB)
                // Highest addr_i = Wrap_Boundary + (Burst_Length x Number_Bytes)
                if (!(&log2_len) &&
                        (((wrap_boundary_o & 12'hfff) + ((burst_length_i + 1) << n_bytes_i)) < (1'b1 << 12))) begin
                    allow_request_o  = 1'b1;     // Allow transaction
                end
                // Boundary violation
                else begin
                    bound_violation_o = 1'b1;
                end

            end

            // BURST_INCR: The final address is Start Addr + Burst_Length x Number_Bytes
            axi_pkg::BURST_INCR: begin
                // check if burst is within 4K range
                if (((addr_i & 12'hfff) + ((burst_length_i + 1) << n_bytes_i)) < (1'b1 << 12)) begin
                    allow_request_o  = 1'b1;     // Allow transaction
                end

                // Boundary violation
                else begin
                    bound_violation_o = 1'b1;
                end
            end

            default:;
        endcase
    end
end

endmodule

/* verilator lint_on WIDTH */
