// Global include file for register interface
// Created for particular use in development process
//

`include "register_interface/typedef.svh"
`include "axi/typedef.svh"

`ifndef GLOBAL_TYPEDEF_SVH
`define GLOBAL_TYPEDEF_SVH

`endif
